module test (
    input [39:0]X,                 // Входная шина X с 40 разрядами (4 группы по 10 разрядов)
	 input [1:0]A,                  // Селектор
    output [9:0]Y);    				  // Выход Y (10 разрядов) для одной группы
	 wire [39:0]TempY;			     // Temp - это просто название переменной, здесь с помощью wire мы просто создали путь шины от входов к выходу
	 assign TempY = X >> A*10;      // Описание работы сдвига. A у нас либо 1, либо 0, но мы добавили умножение на 10, потому как группируем разряды по 10 штук
    assign Y = TempY[9:0];         // [9:0] - позволяет нам выбирать группу разрядов от X0 до X9. То есть выбираем не младший бит, а сразу 10
endmodule                          // Теперь когда A=1, то оно умножается на 10 и двигает группу из 10 разрядов.
