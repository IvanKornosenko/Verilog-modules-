module test (
    input [1:0]X,              // Входная шина X с двумя разрядами
	 input A,                   // Селектор
    output Y);    				 // Выход
	 wire [1:0]TempY;			    // Temp - это просто название переменной, здесь с помощью wire мы просто создали путь шины от входов к выходу
	 assign TempY = X >> A;     // Описание работы сдвига. Мы приваиваем Y значение, полученное при сдвиге. А может быть 1 или 0. 0 - сдвига нет. 1 - сдвиг на 1
    assign Y = TempY[0];       // [0] - означает младший бит (LSB). [1]-старший бит (MSB). В нашем случае мы ориентируемся на младший бит при сдвиге. 
endmodule                      /* По сути, когда A=1, а у нас подано значение 10 (X1X0), то крайний 0 отваливается и мы получаем смещение, в итоге результат 01. 
                                  X1 при смещении сдвигается на позицию X0. В общем такая логика работы у сдвигового MUX*/