module test (input [7:0]X, input [1:0]A, output [1:0]Y);
    MX MX(.Y(Y), .A(A), .X(X));
endmodule
module MX (input [7:0]X, input [1:0]A, output [1:0]Y);
    wire [7:0]Temp = X >> A*2;
    assign Y = Temp[1:0];
endmodule
/* Это наш обычный сдвиговый MUX, который имеет 1 двухразрядный адресный вход и шину X на 8 бит, которая формируется в 4 групы по 2 бита, так как адресный вход двухразрядный. 
Все ничего, но для того, чтобы использовать MUX с другими параметрами, нам придется делать следующее: */

module test (input [7:0]X, input [1:0]A, output [1:0]Y);
    MX1 MX(.Y(Y), .A(A), .X(X));
    MX2 MX(.Y(Y), .A(A), .X(X)); //Добавляем это
endmodule
module MX1 (input [7:0]X, input [1:0]A, output [1:0]Y);
    wire [7:0]Temp = X >> A*2;
    assign Y = Temp[1:0];
endmodule
module MX2 (input [7:0]X, input [1:0]A, output [1:0]Y); //Пишем другой модуль с новыми параметрами и так и будем создавать MX1, MX2,MX3 с разными параметрами
    wire [7:0]Temp = X >> A*2;
    assign Y = Temp[1:0];
endmodule
/* Но наша задача сделать параметризируемый MUX, чтобы не заниматься фигней, которую я описал выше.
   По сути создадим универсальный мультиплексор */

module test (input [3:0]X, input [1:0]A, output Y); // 4-х битная шина X. Адресный вход на 2 бита
    MX #(2) MX(.Y(Y), .A(A), .X(X)); //MX #(2) вот так нужно писать параметры. Это у нас верхний модуль.
endmodule
module MX # (parameter N=2) (input [3:0]X, input [N-1:0]A, output Y); /*      #(parameter N = ) это константа применяемая с появления Verilog 2001. 
                                                                              Она и позволяет сделать нам универсальный MUX, но она будет применяться только в случае,
                                                                              если мы в верхнем модуле не задали параметр. То, что в верхнем модуле - важнее*/
    wire [3:0]Temp = X >> A;
    assign Y = Temp[0];
endmodule
/* Мы создали универсальный MUX с одним параметризируемым адресным входом (A) и с 4-х разрядной шиной (X). С помощью параметра мы задали разрядность 
   адресного входа (A). В общем что бы ни было написано в "MX # (parameter N=2)", parameter будет равен тому, что задали в верхнем модуле ""MX #(2)".  
   Если же в верхнем ничего не задали, тогда выполнится строка "MX # (parameter N=2)"  (Цифра 2 здесь взята просто как пример). */



/*Дальше попробуем сделать MUX еще более гибким, попробуем параметризировать вход "X". */

module test (input [3:0]X, input [1:0]A, output Y); 
    MX #(2) MX(.Y(Y), .A(A), .X(X)); 
endmodule
module MX # (parameter N=2) (input [2**N-1:0]X, input [N-1:0]A, output Y); /* [2**N:0]X. В этом выражении 2**N означает, что мы возводим в степень "N".
                                                                              Но нам нужна шина 4-х разрядная, поэтому делаем (2**N-1), чтобы получилось [3:0] */
    wire [2**N-1:0]Temp = X >> A;
    assign Y = Temp[0];
endmodule



/* Попробуем сделать на большее число разрядов */
module test (input [15:0]X, input [3:0]A, output Y); 
    MX #(4) MX(.Y(Y), .A(A), .X(X)); 
endmodule
module MX # (parameter N=4) (input [2**N-1:0]X, input [N-1:0]A, output Y); // здесь получаем MUX с X шиной на 16 бит и селектор на 3 разряда
    wire [2**N-1:0]Temp = X >> A;
    assign Y = Temp[0];
endmodule



// А теперь добавим еще один параметр "B", который будет влиять на число информационных входов
module test (input [15:0]X, input [3:0]A, output Y); //Если B делаем больше 1, то на наш выход Y тоже будет идти большая разрядность. При B=2, у нас будет [B-1:0]Y
    MX #(.N(4), .B(1)) MX(.Y(Y), .A(A), .X(X));  // MX #(.N(4), .B(1)) Это присваивание параметру N значения 4, а параметру B значения 1
endmodule
module MX # (parameter N=4, B=2) (input [(2**N)*B-1:0]X, input [N-1:0]A, output Y); 
    wire [(2**N)*B-1:0]Temp = X >> A*B; // Сдвиг производим уже группой по 2 (A*B). 
    assign Y = Temp[B-1:0];             
endmodule



//Теперь по сути мы получили универсальный код MUX, их можно размножать и делать какие угодно варианты

module test (input [15:0]X, input [3:0]A, output Y); //то само собой нужно подстраивать под наши новые вводные
    MX #(.N(4), .B(1)) MX(.Y(Y), .A(A), .X(X));
    MX #(.N(2), .B(2)) MX(.Y(Y), .A(A), .X(X));  //Это пример другого MUX с другими параметрами
    MX #(.N(8), .B(4)) MX(.Y(Y), .A(A), .X(X));  //Это пример другого MUX с другими параметрами
endmodule
module MX # (parameter N=4, B=1) (input [(2**N)*B-1:0]X, input [N-1:0]A, output Y); 
    wire [(2**N)*B-1:0]Temp = X >> A*B; 
    assign Y = Temp[B-1:0];             
endmodule



//Рассматриваем дальше то, что мы можем применять. К примеру мы можем применить "localparam"
module test (input [15:0]X, input [3:0]A, output Y); 
    MX #(.N(4), .B(1)) MX(.Y(Y), .A(A), .X(X));
endmodule
module MX # (parameter N=4, B=1) (input [(2**N)*B-1:0]X, input [N-1:0]A, output Y); 
    localparam M = N;                            /*Это тот самый localparam, его можно применять только внутри модуля. Его нельзя изменить извне
                                                   из верхнего модуля. Он привязан  своему модулю, в котором его прописали. Это необходимо для
                                                   того, к примеру, чтобы случайно не накосячить при изменениях параметров в верхнем модуле. */
    wire [(2**N)*B-1:0]Temp = X >> A*B; 
    assign Y = Temp[B-1:0];             
endmodule
  
